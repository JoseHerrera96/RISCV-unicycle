// This file contains the testbench for the Processor module

`timescale 1ns / 1ps

module processor_test;

  // Testbench code goes here

endmodule